LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Adder is

	PORT(x1, x2 : IN STD_LOGIC_VECTOR(3 downto 0);
		  result: OUT STD_LOGIC_VECTOR(3 downto 0);
		  carry : OUT STD_LOGIC_VECTOR);
		  
end Example1


ARCHITECTURE bev of Adder
BEGIN 
	--TODO
END bev;